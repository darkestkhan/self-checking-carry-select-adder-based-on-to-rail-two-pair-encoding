library IEEE;
use IEEE.Std_Logic_1164.all;

entity Half_Adder
is

  port (A, B: in Std_Logic;
        Sum, Carry_Out: out Std_Logic);

end Half_Adder;

architecture Half_Adder_Behav of Half_Adder
is
begin

  Sum <= A xor B;
  Carry_Out <= A and B;

end Half_Adder_Behav;
